module debounce 
    (
        clk,
        in,
        out,
        rst
    );

    input clk;
    input in;
    input rst;

    output reg out;

    always @(posedge clk) begin
    
    end



endmodule
