module twocomplement 
    (
        op1,
        op2,
        out,
    );

    input op1;
    input op2;

    output reg out;

    always @(op1, op2) begin
    
    end



endmodule
